library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ssd_greaterThanComparator is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           X : out  STD_LOGIC);
end ssd_greaterThanComparator;

architecture Behavioral of ssd_greaterThanComparator is

begin


end Behavioral;

