`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:09:25 04/09/2018 
// Design Name: 
// Module Name:    CONTROLLER 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CONTROLLER(
    input CLK,
    input RST,
    input PUSH,
    input POP,
    input [7:0] NUM_IN,
    output [7:0] NUM_OUT,
    output [3:0] SSD_EN,
    output [7:0] EMPTY,
    output [7:0] FULL,
    output [7:0] ST_OV
    );


endmodule
